class minmax_test extends random_test;
    `uvm_component_utils(minmax_test)

function new (string name, uvm_component parent);
    super.new(name,parent);
endfunction : new

    function void build_phase(uvm_phase phase);
        
        super.build_phase(phase);

        // set the factory to produce a add_tester whenever it would produce
        // a random_tester
        command_transaction::type_id::set_type_override(minmax_transaction::get_type());

    endfunction : build_phase
    
endclass