virtual class shape;
	real width;
	real height;
	
	pure virtual function real get_area();
	
	pure virtual function void print();
	
endclass